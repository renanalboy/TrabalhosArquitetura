library verilog;
use verilog.vl_types.all;
entity t_swap is
end t_swap;
